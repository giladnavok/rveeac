
module apb_slave # (
	INIT_FILENAME = "",
	SET_INDEX = 1'b0
) (
	input logic clk,
	input logic rst_n,
	apb_if.slave apb,
	output logic [31:0] mem_o [63:0]
);

logic [31:0] mem [63:0];
assign mem_o = mem;

initial begin
	if (INIT_FILENAME != "") begin
		$readmemh(INIT_FILENAME, mem);
	end 
end

assign apb.rdata = (apb.sel && apb.enable && apb.write == 1'b0) ? mem[(apb.addr/4) % 64] : 32'bx;
assign apb.ready = (apb.sel && apb.enable);
assign apb.slverr = 1'b0;

always_ff @(posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		if (INIT_FILENAME == "") begin
			if (SET_INDEX) begin
				for (int i = 0; i < 64; i++) begin
					mem[i] = i + 32'hffff0000;
				end
			end else begin
				for (int i = 0; i < 64; i++) begin
					mem[i] = '0;
				end
			end
		end
	end else begin
		if (apb.sel && !apb.enable) begin
			if (apb.write) begin
				case (apb.strb) 
					4'b1111: mem[apb.addr/4] <= apb.wdata;
					4'b0011: mem[apb.addr/4][15:0] <= apb.wdata[15:0];
					4'b0001: mem[apb.addr/4][7:0] <= apb.wdata[7:0];
					default: mem[apb.addr/4] <= apb.wdata;
				endcase
			end
		end
	end
end
endmodule
