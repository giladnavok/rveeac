
module controller (


);
