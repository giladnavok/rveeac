
module tbFetchUnit;

// IMEM interface
logic clk;
logic resetN;
logic [7:0] addr;
logic write;
logic [31:0] din;
logic [31:0] dout;

MemorySubmodule 
imem (

endmodule
